library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity VGA_RETO is
    port(
        CLK : in std_logic; B0, B1, B2, B3, B4, B5, B6, B7, B8, B9 : in std_logic_vector(7 downto 0);
        R, G, B : out std_logic_vector(3 downto 0); 
        VS, HS : out std_logic
    );
end VGA_RETO;

architecture behav of VGA_RETO is

    component DIVISOR_CLOCK is
        generic( pulsos : integer := 1);
        port(clk_in: in std_logic; clk_out : out std_logic);
    end component;

    signal clk_25M : std_logic;
    signal HS_signal, VS_signal, flag_hs, flag_vs, flag_check : std_logic;
    signal R_temp, G_temp, B_temp : std_logic_vector(3 downto 0);
    signal spox : std_logic_vector(9 downto 0);
    signal spoy : std_logic_vector(8 downto 0);

 
    constant DIGIT_WIDTH : integer := 60;  -- Ancho de cada número
    constant DIGIT_HEIGHT : integer := 60; -- Alto de cada número
    constant DIGIT_SPACING : integer := 0; 
    constant START_X : integer := 20;      -- Posición inicial en X
    constant START_Y : integer := 100;     -- Posición inicial en Y
	 constant START_X_BARRA : integer := 20; 
	 constant START_Y_BARRA : integer := 170;
	 constant BAR_WIDTH : integer := 0;

    type digit_0_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_0 : digit_0_array := (
		 
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		
	);

	type digit_1_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_1 : digit_1_array := (
		 
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000111100000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000111111000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
	
	);

	type digit_2_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_2 : digit_2_array := (
		
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000011000000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000111110000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		 
	);

	type digit_3_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_3 : digit_3_array := (
		 
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		 
	);

	type digit_4_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_4 : digit_4_array := (
		
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000001110000000000000000000000000000",
		 "000000000000000000000000000010110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000111111000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
	);

	type digit_5_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_5 : digit_5_array := (
		 
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000111110000000000000000000000000000",
		 "000000000000000000000000000110000000000000000000000000000000",
		 "000000000000000000000000000111100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000100110000000000000000000000000000",
		 "000000000000000000000000000111100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		 
	);

	type digit_6_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_6 : digit_6_array := (
		 
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110000000000000000000000000000000",
		 "000000000000000000000000000111100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		 
	);

	type digit_7_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_7 : digit_7_array := (
		
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000111110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000001100000000000000000000000000000",
		 "000000000000000000000000000011000000000000000000000000000000",
		 "000000000000000000000000000011000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		 
	);

	type digit_8_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_8 : digit_8_array := (
		
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		
	);

	type digit_9_array is array (0 to 59) of std_logic_vector(59 downto 0);
	constant digit_9 : digit_9_array := (
		
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011110000000000000000000000000000",
		 "000000000000000000000000000000110000000000000000000000000000",
		 "000000000000000000000000000110110000000000000000000000000000",
		 "000000000000000000000000000011100000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--20
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",--10
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000"
		
	);

	type bar_0_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_0 : bar_0_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000"
	);
	
	type bar_1_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_1 : bar_1_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );


	
	type bar_2_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_2 : bar_2_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );

	
	type bar_3_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_3 : bar_3_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );
	
	type bar_4_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_4 : bar_4_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );

	
	type bar_5_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_5 : bar_5_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );

	
	type bar_6_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_6 : bar_6_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );


	
	type bar_7_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_7 : bar_7_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );

	
	type bar_8_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_8 : bar_8_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );

	
	type bar_9_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_9 : bar_9_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 );
		 
		 
	type bar_10_array is array (0 to 249) of std_logic_vector(59 downto 0);
	constant barra_10 : bar_10_array := (
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",
		 "000000000000000000000000000000000000000000000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001100000000000000001100000000000000000000",---
		 
		 "000000000000000000001100000000000000001100000000000000000000",---
		 "000000000000000000001101111111111111101100000000000000000000",--
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001101111111111111101100000000000000000000",
		 "000000000000000000001100000000000000001100000000000000000000",
		 "000000000000000000001111111111111111111100000000000000000000",--
		 "000000000000000000001111111111111111111100000000000000000000"---
		 
		 
	);




begin

		U0: DIVISOR_CLOCK port map (CLK, clk_25M);
		flag_check <= flag_vs and flag_hs; -- comprobamos que estamos en el display time de HS y VS

    process (clk_25M)
        variable x, y, i : integer;
        variable pixel_on : std_logic;
		  variable local_x, local_y : integer;
		  variable local_x_bar, local_y_bar : integer;
    begin
        if rising_edge(clk_25M) then
            x := to_integer(unsigned(spox));
            y := to_integer(unsigned(spoy));

            R_temp <= "0000";
            G_temp <= "0000";
            B_temp <= "0000";
            
            -- Recorrer los 10 números
            for i in 0 to 9 loop
                if (x >= START_X + i * (DIGIT_WIDTH + DIGIT_SPACING)) and 
                   (x < START_X + i * (DIGIT_WIDTH + DIGIT_SPACING) + DIGIT_WIDTH) and 
                   (y >= START_Y and y < START_Y + DIGIT_HEIGHT) then
                    
                    -- Obtener la posición dentro del número
                    local_x := x - (START_X + i * (DIGIT_WIDTH + DIGIT_SPACING));
                    local_y := y - START_Y;

                    case i is
                        when 0 => pixel_on := digit_0(local_y)(59 - local_x);
                        when 1 => pixel_on := digit_1(local_y)(59 - local_x);
                        when 2 => pixel_on := digit_2(local_y)(59 - local_x);
                        when 3 => pixel_on := digit_3(local_y)(59 - local_x);
                        when 4 => pixel_on := digit_4(local_y)(59 - local_x);
                        when 5 => pixel_on := digit_5(local_y)(59 - local_x);
                        when 6 => pixel_on := digit_6(local_y)(59 - local_x);
                        when 7 => pixel_on := digit_7(local_y)(59 - local_x);
                        when 8 => pixel_on := digit_8(local_y)(59 - local_x);
                        when 9 => pixel_on := digit_9(local_y)(59 - local_x);
                        when others => pixel_on := '0';
                    end case;

                    
                    if pixel_on = '1' then
                        R_temp <= "1111";
                        G_temp <= "1111";
                        B_temp <= "1111";
                    end if;
                end if;
            end loop;
				
				for i in 0 to 9 loop
					if ( x >= START_X + i * (DIGIT_WIDTH + DIGIT_SPACING)) and 
                   (x < START_X + i * (DIGIT_WIDTH + DIGIT_SPACING) + DIGIT_WIDTH) and 
						 (y > START_Y_BARRA and y < 420) then
						 
						local_x := x - (START_X_BARRA + i * (DIGIT_WIDTH + DIGIT_SPACING));
                  local_y := y - 170;
						
						case i is
                        when 0 => 
									case b0 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
									
                        when 1 => 
									case b1 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 2 => 
									case b2 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 3 => 
									case b3 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 4 => 
									case b4 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 5 => 
									case b5 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 6 => 
									case b6 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 7 => 
									case b7 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 8 => 
									case b8 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when 9 => 
									case b9 is
										when "00110000" => pixel_on := barra_0(local_y)(59 - local_x);
										when "00110001" => pixel_on := barra_1(local_y)(59 - local_x);
										when "00110010" => pixel_on := barra_2(local_y)(59 - local_x);
										when "00110011" => pixel_on := barra_3(local_y)(59 - local_x);
										when "00110100" => pixel_on := barra_4(local_y)(59 - local_x);
										when "00110101" => pixel_on := barra_5(local_y)(59 - local_x);
										when "00110110" => pixel_on := barra_6(local_y)(59 - local_x);
										when "00110111" => pixel_on := barra_7(local_y)(59 - local_x);
										when "00111000" => pixel_on := barra_8(local_y)(59 - local_x);
										when "00111001" => pixel_on := barra_9(local_y)(59 - local_x);
										when "00111010" => pixel_on := barra_10(local_y)(59 - local_x);
										when others => pixel_on := barra_0(local_y)(59 - local_x);
									end case;
                        when others => pixel_on := '0';
                    end case;
						  -- Si el bit está activo, pintar en blanco
                    if pixel_on = '1' then
                        R_temp <= "1111";
                        G_temp <= "1111";
                        B_temp <= "1111";
                    end if;

					 end if;
				end loop;
				
				
        end if;
    end process;
	 
	 
		--      _:HS SIGNAL:_
		-- Pulse width : 0-95
		-- back porch : 95-143
		-- display time : 143 - 783
		-- front porch : 783 - 799 pulsos 
		P0 : process(clk_25M)
			variable contador_hs : integer := 0;
			variable posicion_x : integer := 0;
			begin
				if rising_edge (clk_25M) then
					contador_hs := contador_hs + 1;
					if contador_hs < 96 then -- pulse width
						HS_signal <= '0';
						flag_hs <= '0';
					elsif contador_hs < 144 then  -- back porch
						HS_signal <= '1';
						flag_hs <= '0';
					elsif contador_hs < 784 then  -- display time
						HS_signal <= '1';
						flag_hs <= '1';
						posicion_x := posicion_x +1;
					elsif contador_hs < 800 then  -- front porch
						HS_signal <= '1';
						flag_hs <= '0';
					else
						contador_hs := 0;
						HS_signal <= '0';
						flag_hs <= '0';
						posicion_x := 0;
					end if;
				else
					contador_hs := contador_hs;
				end if;
				
				spox <= std_logic_vector(to_unsigned(posicion_x,10));
		end process;
		
		HS <= HS_signal;
		
		
		
		
		--      _:VS SIGNAL:_
		-- Pulse width : 0-1
		-- back porch : 1-30
		-- display time : 30 - 510
		-- front porch : 510 - 520 líneas de VS 
		P1 : process(HS_signal) 
			variable contador_vs : integer := 0;
			variable posicion_y : integer := 0;
			begin
				if falling_edge (HS_signal) then -- es falling edge porque en falling_edge de HS, VS empieza
					contador_vs := contador_vs +1;
					if contador_vs < 2 then
						VS_signal <= '0';
						flag_vs <= '0';
					elsif contador_vs < 31 then
						VS_signal <= '1';
						flag_vs <= '0';
					elsif contador_vs < 511 then
						VS_signal <= '1';
						flag_vs <= '1';
						posicion_y := posicion_y +1;
					elsif contador_vs < 521 then
						VS_signal <= '1';
						flag_vs <= '0';
					else
					contador_vs := 0;
						VS_signal <= '0';
						flag_vs <= '0';
						posicion_y := 0;
					end if;
				else
					contador_vs := contador_vs;
				end if;
				spoy <= std_logic_vector(to_unsigned(posicion_y,9));
		end process;
		
		VS <= vs_signal;
		

    -- Asignación de las señales de salida
    R <= R_temp;
    G <= G_temp;
    B <= B_temp;
    HS <= HS_signal;
    VS <= VS_signal;
	 
	 

end behav;
